// SPDX-License-Identifier: SHL-2.1

module clarigggz_core (
    input wire clk,
    input wire rst_n,
    // RISC-V signals
    output wire [63:0] pc,
    input wire [31:0] instruction
);

    // Placeholder for custom RISC-V RV64GCV implementation
    
endmodule
